module baud_gen
  import definitions_pkg::*;
  ( 
    input   logic clk, 
    input   logic rstN,
    output  logic baud_tick
  );  

  

endmodule: baud_gen