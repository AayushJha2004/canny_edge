module sqrt_22b (
    input  logic [21:0] value,     
    output logic [10:0] sqrt    
);
    
endmodule
