module gaussian_filter
  import definitions_pkg::*;
(
  
);
endmodule: gaussian_filter